module CONFF (
    input [31:0] IR,
    output reg [31:0] to_Control 
);

reg [4:0] C2,
