module bus()
    wire[31:0] input_wire
    wire[4:0] output_wire
    input_wire[0] = R0out
    
    encoder_32_5 encoder()
endmodule