include "./reg_test.v"
module bus;

endmodule;