module bus(
    encoder_32_5 A();
    
    reg_32bit R0(clk,clear,r0_enable,buscontents,r0_out);
    
    
    32_1_decoder B();

)
endmodule
module datapath(

)
end datapath