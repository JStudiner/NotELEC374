module ELEC374ProjectSim(
    input wire A,
    output reg B
);
endmodule