module 32_1_decoder();
endmodule;